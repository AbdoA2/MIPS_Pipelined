import cache_def::*;
module ICache(input logic clk, reset,
              input cpu_req_typeI cpu_req,
              output cpu_result_type cpu_result,
              output mem_req_typeI mem_req,
              input mem_result_type data);
  
  cache_data_type rd1, rd2;
  cache_req_type d_req1, d_req2, t_req1, t_req2;
  tag_type wt, rt1, rt2;
  logic[1:0] offset;
  logic[31:0] instr;
  
  assign offset = cpu_req.addr[3:2];
  
  data_mem way1(clk, reset, d_req1, mem_result.data, rd1);
  data_mem way2(clk, reset, d_req2, mem_result.data, rd2);
  
  tag_mem tag1(clk, reset, t_req1, wt, rt1);
  tag_mem tag2(clk, reset, t_req2, wt, rt2);
  
  
  typedef enum logic {idle, fetch} state_type;
  state_type state, nextstate;
  
  // read data
  assign data1 = offset[1]? (offset[0]? rd1[127:96] : rd1[95:64]) : (offset[0]? rd1[63:32] : rd1[31:0]);
  assign data2 = offset[1]? (offset[0]? rd2[127:96] : rd2[95:64]) : (offset[0]? rd2[63:32] : rd2[31:0]);
  
  // check hit
  assign h1 = (rt1.tag == cpu_req.addr[31:8] & rt1.valid);
  assign h2 = (rt2.tag == cpu_req.addr[31:8] & rt2.valid);
  assign hit = h1 | h2;
  
  // choose the instruction
  assign instr = h1? data1 : data2;
  
  always_comb begin
    
    // default values write enable must be zero and assign the cpu requested address
    d_req1 <= {cpu_req.addr[7:4], 1'b0};
    d_req2 <= {cpu_req.addr[7:4], 1'b0};
    t_req1 <= {cpu_req.addr[7:4], 1'b0};
    t_req2 <= {cpu_req.addr[7:4], 1'b0};
        
    if (state == idle) begin
      if (cpu_req.valid == 1'b1) begin
        
        if (hit) begin
          
          cpu_result.data <= instr;
          cpu_result.ready <= 1'b1;
          mem_req.valid <= 1'b0;
          nextstate <= idle;
          
        end
        else begin
          
          cpu_result.ready <= 1'b0;
          mem_req.addr <= {cpu_req.addr[31:4], 4'b0};
          mem_req.valid <= 1'b1;
          nextstate <= fetch;
          
        end
      end
    end
    else begin
      if (mem_result.ready) begin
        if (rt1.valid == 1'b0) begin
          d_req1.we <= 1'b1;
          rt1.dirty <= 1;
          rt2.dirty <= 0;
        end
        else if (rt2.valid == 1'b0) begin
          d_req2.we <= 1'b1;
          rt2.dirty <= 1;
          rt1.dirty <= 0;
        end
        else if (rt1.dirty) begin
          d_req2.we <= 1'b1;
          rt2.dirty <= 1;
          rt1.dirty <= 0;
        end
        else begin
          d_req1.we <= 1'b1;
          rt1.dirty <= 1;
          rt2.dirty <= 0;
        end
        
        cpu_result.ready <= 1'b1;
        mem_result.valid <= 1'b0;
        nextstate <= idle;
      end
      else begin
        nextstate <= fetch;
      end
    end
  end
  
  always_ff @ (posedge clk) begin
    if (reset) state <= idle;
    else state <= nextstate;
  end
  
  
endmodule
